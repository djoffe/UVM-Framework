//----------------------------------------------------------------------
//   Copyright 2013 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//                   Mentor Graphics Inc
//----------------------------------------------------------------------
// Project         : gpio interface agent
// Unit            : Sequence library
// File            : gpio_random_sequence.svh
//----------------------------------------------------------------------
// Creation Date   : 05.12.2011
//----------------------------------------------------------------------
// Description: This sequence exists to support the python based test
//    bench generator.  The test bench generator instantiates a random
//    sequence for each ACTIVE agent added to the bench.
//
//----------------------------------------------------------------------
//
class gpio_random_sequence #(int READ_PORT_WIDTH=4, int WRITE_PORT_WIDTH=4) extends 
    gpio_sequence_base #( READ_PORT_WIDTH, WRITE_PORT_WIDTH );

  `uvm_object_param_utils( gpio_random_sequence #(READ_PORT_WIDTH, WRITE_PORT_WIDTH))

// ****************************************************************************
  function new( string name ="");
    super.new( name );
  endfunction

// ****************************************************************************
  task body();
     `uvm_info("SEQ","REPLACE GPIO_RANDOM_SEQUENCE WITH YOUR EXTENSION OF GPIO_SEQUENCE",UVM_NONE);
  endtask

endclass
