
import uvm_pkg::*;
import qvip_usb3_pipe_example_bench_test_pkg::*;

module hvl_top;


initial run_test();

endmodule

