/*****************************************************************************
 *
 * Copyright 2007-2015 Mentor Graphics Corporation
 * All Rights Reserved.
 *
 * THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY INFORMATION WHICH IS THE PROPERTY OF 
 * MENTOR GRAPHICS CORPORATION OR ITS LICENSORS AND IS SUBJECT TO LICENSE TERMS.
 *
 *****************************************************************************/


module ethernet_dummy_dut (
                        reset,
                        clk_0,
                        txd,
                        txc,
                        clk_1,
                        rxd,
                        rxc
                        );
  import uvm_pkg::*;
  import mvc_pkg::*;
  import mgc_ethernet_v1_0_pkg::*;
 
   input         reset;
   input         clk_0;
   output [31:0] txd;
   output [3:0]  txc;
   input         clk_1;
   input [31:0]  rxd;
   input [3:0]   rxc;
    
   parameter ERRONEOUS_FRAMES_ON = 0;
   parameter EEE_ENABLED = 0;
   
   reg [31:0]    txd;
   reg [3:0]     txc;
   
   initial
     begin
        txd = 32'h07070707;
        txc = 4'hF;
        repeat (11) @(clk_0);
        
        if(ERRONEOUS_FRAMES_ON)
        begin
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h1acfd5fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h65878651;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hff000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000ffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10100000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10101010;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10101010;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10101010;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10101010;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10101010;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10101010;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10101010;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10101010;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10101010;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10101010;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h36871010;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fdb017;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h97d555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'haa9d4e73;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000029;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00ffffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0b0b0b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0b0b0b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0b0b0b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0b0b0b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0b0b0b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0b0b0b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0b0b0b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0b0b0b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0b0b0b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0b0b0b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf1b0b0b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfdb35474;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'hd55555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h7125100c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000030a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hadf30081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e3e3e3e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e3e3e3e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e3e3e3e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e3e3e3e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e3e3e3e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e3e3e3e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e3e3e3e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e3e3e3e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e3e3e3e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e3e3e3e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e3e3e3e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf3709bbe;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h8b4a95d5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00361e3a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffff0000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h580081ff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000000d1;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h09090900;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h09090909;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h09090909;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h09090909;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h09090909;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h09090909;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h09090909;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h09090909;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h09090909;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h09090909;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h09090909;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb954d709;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0707fd18;
          txc <= 4'he;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h52d5d555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he93f65e3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hff000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000ffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f1f0000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f1f1f1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f1f1f1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f1f1f1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f1f1f1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f1f1f1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f1f1f1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f1f1f1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f1f1f1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f1f1f1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f1f1f1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfcc41f1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fd0497;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h71d55555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb53faf6b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000007b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h81ffffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00d5dc00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h90505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfda066a4;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hc8d55555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4321ad08;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000000db;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00ffffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h44505050;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfd1b3a4f;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h512e1cd5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00fde223;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffff0000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc20081ff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000053;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16161600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16161616;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16161616;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16161616;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16161616;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16161616;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16161616;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16161616;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16161616;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16161616;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16161616;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6d83ed16;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0707fddd;
          txc <= 4'he;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha9a6d555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h175b6e68;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hff000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0081ffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00002b37;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95950000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf4709595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fd8834;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h08d55555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6988a4c0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000000c7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00ffffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hba000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbabababa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbabababa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbabababa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbabababa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbabababa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbabababa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbabababa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbabababa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbabababa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbabababa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h52bababa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfd2acf5a;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h861e8ebd;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000b0b2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd6bc0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3155effe;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf54d2ed5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h004b4e05;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffff0000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000000ff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a9a9a00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a9a9a9a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a9a9a9a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a9a9a9a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a9a9a9a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a9a9a9a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a9a9a9a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a9a9a9a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a9a9a9a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a9a9a9a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a9a9a9a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0c73bf9a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0707fd26;
          txc <= 4'he;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1feed555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5e58ff62;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hff000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000ffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdede0000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdededede;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdededede;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdededede;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdededede;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdededede;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdededede;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdededede;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdededede;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdededede;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdededede;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h85f4dede;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fd9ab5;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h61d55555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h327d0a63;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000060;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00ffffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46464646;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46464646;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46464646;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46464646;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46464646;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46464646;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46464646;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46464646;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46464646;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46464646;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h40464646;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfd5c18c9;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haa8d0432;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000c82b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9aad0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4dc536d4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h83bd118b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000b375;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43434343;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd2e05946;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h5555fb07;
          txc <= 4'h3;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h11e852d5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h003ea7d0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffff0000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc50081ff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000000d1;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5d5d5d00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5d5d5d5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5d5d5d5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5d5d5d5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5d5d5d5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5d5d5d5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5d5d5d5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5d5d5d5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5d5d5d5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5d5d5d5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5d5d5d5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3af69b5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0707fd66;
          txc <= 4'he;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h55fb0707;
          txc <= 4'h7;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h605cd555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h365249ea;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hff000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000ffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haeae0000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haeaeaeae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haeaeaeae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haeaeaeae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haeaeaeae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haeaeaeae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haeaeaeae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haeaeaeae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haeaeaeae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haeaeaeae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haeaeaeae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h49d1aeae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fd4c92;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'hfb070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8cd55555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h34845834;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000000bb;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h81ffffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00185f00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h01959595;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfddc2373;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hcf85190f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00002ca6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he5bc0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h54545454;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h54545454;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h54545454;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h54545454;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h54545454;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h54545454;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h54545454;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h54545454;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h54545454;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h54545454;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h54545454;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd698ee68;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h842b190d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000541b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b9b9b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b9b9b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b9b9b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b9b9b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b9b9b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b9b9b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b9b9b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b9b9b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b9b9b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b9b9b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b9b9b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b9b9b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfce87505;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb6487c17;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000063f2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hecececec;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hecececec;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hecececec;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hecececec;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hecececec;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hecececec;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1c17ecec;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fd5985;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha679b0cc;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000a866;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5f000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfdf191a8;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h8001d5fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h010000c2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hff000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0081ffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h08884a4f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h52e00100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h20e00000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fd1464;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'hdfd555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hf3e96b2f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000001e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h88ffffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc3100008;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00405268;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h15000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfd7a8d36;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'hd55555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h00c28001;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h01000888;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00006cd4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha38d3b5b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hffdf53d5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00df9ced;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffff0000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he30081ff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0008888b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h56297410;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000000b2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1719c200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0707fd97;
          txc <= 4'he;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hf8f6d555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h35f606d0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hff000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0081ffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h088889de;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hddb91000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000fc7c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc6b10000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fd7364;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h01d55555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000c280;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000001;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h88ffffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h96010008;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000000d3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfd53bd45;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h09d55555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6e884d77;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000002;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h81ffffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h88fcbb00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf2100008;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h001d7038;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hee000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfde4305f;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc28001d5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00010000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffff0000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf90081ff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000888b1;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h003c3901;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h03640a00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0707fd97;
          txc <= 4'he;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8001d555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h010000c2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hff000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0888ffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h66410100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46e20000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fdfb0f;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h01d55555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000c280;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000001;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h81ffffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h88d12e00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h84010008;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000077;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdc000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfd7199bc;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00c28001;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h01000888;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000fdef;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h60136b72;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc28001d5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00010000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffff0000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd20081ff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000888ab;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00712201;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc06aaa00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0707fdb1;
          txc <= 4'he;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8001d555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h010000c2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hff000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0888ffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha4860100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h65050000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fd720b;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h01d55555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000c280;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000001;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h88ffffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0c010008;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000000ea;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h96000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfdbbb9c7;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00c28001;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h01000888;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00002250;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1cffcdd5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00c28001;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd63a0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h01000888;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000077f2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc4989f5b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h5555fb07;
          txc <= 4'h3;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc28001d5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00010000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffff0000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h230081ff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0008888c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00ae3e01;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb30efa00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0707fd2c;
          txc <= 4'he;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h55fb0707;
          txc <= 4'h7;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8001d555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h010000c2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hff000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0888ffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h27d80100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5b8f0000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fdd8d3;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'hfb070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h55555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf2d55555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h02f09df0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000000c2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h88ffffff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h40100008;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00b21c69;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf8000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfd1687af;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he15675de;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000059ef;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7a6f0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10000888;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h08f779e3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7c6231b5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00c28001;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h01000888;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000c0d3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000c0d3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h38b8c299;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00c28001;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb4b00081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h506b0888;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fd100a;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00c28001;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h01000888;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000c0f4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hab307430;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h956f8718;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00005138;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h20f40081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf9113900;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h29606486;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb5577e2d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc1899027;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4a2cc8aa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h48e5cbbd;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7b1326e0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfaeecc54;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7aa94859;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h74e4d254;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbe2ae7a7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h40c98052;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc058d8f3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h019db884;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h578a138d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfd3f8938;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4d47b704;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000ff2b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0d1d0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd4f83200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h177f4b1a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hced346d9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0e564f11;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbeb374d5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffe58533;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb280d15f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1cb81802;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha6bd808b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h97f405d3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h87642f8a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'had5aae02;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h22ba990c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4603338b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h367618c0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00004afb;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfa4a0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf3c63600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3347b8a0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h64343ead;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc4c31ab3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8cd46f2b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h475115b1;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hce0efb3d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4e810ee0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha0e21af6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7612008a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07574bba;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h45b0db18;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9b2591d4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb2b9ab27;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc20867b3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc1026fa9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00003952;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he1ea3800;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hcda2ca47;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0c18fa98;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10873f40;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf0bbecee;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4ae7ced5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h36b6aea5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h13c2cbc1;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h24c3208e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb7a7f0c9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdcf43f3a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha345089e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h50e50218;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7a7e82eb;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he8ee8ab3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fd2796;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha7f61482;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000f97c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6c2e3200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2a126cb6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h93e71726;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8b746d48;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h31bc7a4d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07dd285a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h268f58bb;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd495de5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5a5ca334;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfd164144;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h68d30159;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h854f1634;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h98ae5c5c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3f218a1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd2584c6f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00009687;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h25463600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8444cb07;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2d1583fb;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc5ab8ebd;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h33f28c88;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h560a545e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf1c8da27;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9e3a898;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf9618501;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hcdc1dd69;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h67cc9a06;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb618b1ef;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6c820a2f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6e5528db;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h94dcd130;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha60d82b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00006af3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf9610081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0b6f3700;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hda508c16;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0595aea9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0a21a5f7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc7177e24;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h28286dfa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd803b3f4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc4de48aa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7c036573;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8e10228a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc548bcaf;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbf1e2a00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4dcb496b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8935ac18;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb866e442;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0707fdc2;
          txc <= 4'he;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f501aa2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00004191;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h52363200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4936a6e4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc5a7a381;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3ca2a774;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb1ae609a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0a4edd6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbc51e21b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hecf1bd3a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd6ddc193;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9ec4490b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h054427d9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h946b4fe9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1a464b06;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h61a74996;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h793e24e9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00009ac2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1b080081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h51ab3600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h87cce17d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h82021300;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7cc4a8b9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hacb445ad;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7ac888b8;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha127f34e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h664c652c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2276adb5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h78f6b8b5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb25b3d85;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf7d8c033;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb9b669b6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1c5d7237;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd7f9233d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc085bc24;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00009b2e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h663c3600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h952df05c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h588d7754;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha5f061e9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha00d5880;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb372efc2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc8832bac;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd306b4f2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h52202ab3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h98ee7e20;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h37e2af8a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfc2b3c55;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h76a6e5dc;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h38d1ed15;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc239c3fc;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he6d23e09;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00005f42;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7e790081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hed0e3200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f4b94e9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3b8d1b91;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5a469cf2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbd6cbc06;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2a5f1a56;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h49fc19f1;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h013fc5f6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7b727716;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h239757f7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he0af3e8f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h45926884;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbfdeaf11;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc6e8d183;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8abf8d0a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000d2ff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2fb43600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9554a744;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1b5924bc;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he4909819;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8a36aa0b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha532dd30;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he060b983;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h404c1bd2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1fecc160;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf5d9cb7f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7a634be3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbd16205a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2108b233;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4f6b4c9d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6055f008;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6604ab49;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000306;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5ca40081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00943500;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h49d3928a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc4f2a0f4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hcdbe6537;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha7654d93;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h95003025;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h89818676;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h37d5ca29;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha3107e14;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h80e1b429;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h811e27ce;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h282e9311;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h22ad31ad;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h410a6f94;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfd77b956;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hed28fc18;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00005e5c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb0a60081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h51643200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he3477cf2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h94d4ff64;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbcdaa8ba;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hecde7073;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h903b51b6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2b14e0ef;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h48fb2a10;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6e319d2a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5da2e3c7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc58b4299;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc62bb2af;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1cf34c29;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf789c2ce;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb5411cde;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00004e38;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf9d03600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h93143d87;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h29827ff9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h27bde451;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdb1d2080;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haf98c3aa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4ae3fca7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1c016776;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h66b8eb7c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h96b41db2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9e7d534f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc4bd6122;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hef7001ad;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h277888ad;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdf293142;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h388ffa09;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00003aec;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hadc33400;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb2d45a75;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb4aea41e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5b53f721;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6d31376b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3f212dbe;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h83fa0db6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1a011d1f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1a49b257;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2e5fbfe2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0598e18c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h595358f6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h099a409f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h874584ef;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fd3297;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h15ce459c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000b9f6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46c33200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7afb4638;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf4c26f54;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4e845dcb;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5e7f9089;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'heeadb8b8;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h30ed0623;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7f72868b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7510fead;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc4a44a5d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h06f69f4b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h855781f2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha5102926;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha2976303;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h29f9acf6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000688d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10f33600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbaa7b4af;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h29da4ea0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7002d5ae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6e334005;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4dcc37d5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he71dda70;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h27439ecf;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbf110cdc;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbf5f0aed;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h09aa2de3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h64fed481;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h97517de1;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd73ca7c0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2662284a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc4b7243f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000e928;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdd2c3300;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5ab07a9a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h68c56ba8;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2f410100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he2f018b1;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7decfc76;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hab7825b8;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha7f7ae71;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'heb50241b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he93f86dc;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h60a823f7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46eb8c39;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1fff0637;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha65ed740;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0707fd85;
          txc <= 4'he;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5d8891be;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000dd75;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h896f3200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h56d0d0e0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4a1b88c0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h026201d2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h252c5d78;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha0ea3d38;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd6be74ce;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'head1b419;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7e34fd9f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h87e5544d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9356f5d9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h37a2b97c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf5d7bbab;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc6f06a5e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc5c269ef;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000051c7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7b300081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h72863600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc4ad5b13;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h88ccc7a6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf1ddce1d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd9c59f5a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4cb1c63e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0c74c7f7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he9adb585;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5fcf79e8;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf4dd1e6a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h62575874;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hef4fc42e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7b59315e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4496de8a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h908b1254;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f0765a4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000b581;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8ffc0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h18583200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h23ddbec9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4e7a8453;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h20c9b371;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hab93c6f9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf5026f06;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8a536d0a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he749c0ff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haca595c0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbcb25fe7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdc5410b1;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc6972907;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h35c53406;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h85dfaf40;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h962a5020;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000775;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7d3c0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h28673200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h65af050f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h513fc6ad;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h775e7f9f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hef08f21c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'head3fcd4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfdafe91e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4a1ef592;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9182ec31;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfba76dcd;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9de779ef;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h041a8d4d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbb153371;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'heef96748;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h065825fb;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000d8b3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h49ac0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h14fb3600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9890ecad;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a9e582f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h73b61356;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h80d554e6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he9a0ae69;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6cfb6ec6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf25b250e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfe75889b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2b176e95;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h03351038;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h48f85405;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdbfaddb0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haac145b8;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he784ab4b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdd998878;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00006718;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h96070081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdc9d3100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfe0994bf;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha38d3e89;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h67ac41eb;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haba3d068;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdc532e89;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16fde707;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5041b5c2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc64ba081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43a5153f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h02ca05a7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9061bdf9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h47a5589b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfd7f1a20;
          txc <= 4'h8;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdb02403b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00005288;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46010081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8e9f3200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hba245922;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h991492b6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07c20380;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7b9ebe4d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc23c1054;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he8866bea;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha1d8455b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h64fb3388;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5bd9c2cc;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5b67fdd6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc8c17d58;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h299be7d7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0c8a0342;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6f72a9bb;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00002cb0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6f520081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb05d3600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd0f9de50;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'had92e5b4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd3a86850;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h46af40f4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb5c1b5af;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0a9bb2c3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hace83ff0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfa11069a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc91dd8f4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4fecee1c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9fffc722;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h816abb17;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd8b7d4ba;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8af15971;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3938b19d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000ee3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h456c3000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h713cb7c1;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h11b2f1a5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9d25bb17;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h565a404e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h18f156e9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb7e558e3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h42f2a1e5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hcc586833;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfbf33612;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h52ca79b0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbf42b797;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9b56a2c5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h07fd8d72;
          txc <= 4'hc;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0d2cf072;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000e56a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h23743200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc5e961dc;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7715f074;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfbf65ed4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha95dfc5c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha2a2f4e3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd631b69b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hacae903b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0d8628cc;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfb9439de;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4ddb5bd9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1eacb734;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h04a278e8;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h469a43bc;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hba5146e4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000a53;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h63823600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16b01519;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0ded8fea;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he5d4365f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5c6e0883;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfdff6cc6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf95b3401;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2be7ecff;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h330a6d1c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h125d413b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf9544734;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3c2e53fb;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h92b74a97;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha6002af6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6f0aeca3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h213f4f7e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00003a1d;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h116e0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb22c2f00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1ce481df;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2461398e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha45cbd1a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he6caf540;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'heb599503;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd1942e83;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h64aa013f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha273c633;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h574e8492;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5a7512ba;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbb9ccf14;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2cc2c09a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0707fd3e;
          txc <= 4'he;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h653d4760;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h000073e3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbb140081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43173200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'haf66b1ab;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h488613ad;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5c678adf;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h165ad324;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7c54f659;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3a225b95;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9a7d9ccc;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f0e8a71;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0b76f794;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h595ca831;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5789013f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6d4aabe5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h711290a7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbecc46db;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00002427;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hfd920081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e043600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc2a2abc3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7bd0c2c9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb209d765;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he1c310f4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h694315de;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4f72a453;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h007c33cf;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0c1e2826;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4cfcac12;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9d2f7694;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6a8aec35;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbb5820c6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4754f228;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd512ceab;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc60ad148;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000f553;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h375d0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h730a2e00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1f0f0b7b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h86a4d4d5;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5b30d0e4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5472ef2f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb7cd0fa7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb2f964f6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hcc4397ae;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6d998a57;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6f573634;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc8440b14;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2ce33a7e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h694c56e6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4690d8e0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000232;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9ecc0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h2e4b3200;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8e510ab6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h77ac901e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h29446e29;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h257970cb;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9ad8a69f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hecac022b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1e09655f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hff05dd9e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h9bfabc51;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43a4e2b1;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hcf2e7eef;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6172260c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5320f9c3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbca58804;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000594f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd8b03600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha8949316;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h45974fbf;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc180c105;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6c1e19c3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5c0ceeaa;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7c41d59c;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3eae202b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'heea1c9e8;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h21ce972e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5be192a1;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h43e2a094;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6e27698f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hed67f610;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8a2bd8f3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd555fe55;
          txc <= 4'h2;
          @ clk_0;
          txd <= 32'hbc4c551b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000670e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h672c0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha0aa3600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hf8774e28;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hd2ea3a32;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hbf7bd084;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he18ca52b;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6eb0e6ca;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h271a1ce4;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hff6729b2;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h585c1457;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h01d63c94;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h79739931;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb811c8cf;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h657f4fa9;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h53666483;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h33a4548e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd555fe55;
          txc <= 4'h2;
          @ clk_0;
          txd <= 32'h00c28001;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000100;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h01000888;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00002948;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hc5e72271;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h5a3c9d67;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000c9ef;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha4d60081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h3e2e3600;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h53faec25;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h45d2861e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'ha7fe172c;
          txc <= 4'h4;
          @ clk_0;
          txd <= 32'h75a89e28;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hdc852d87;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h7b6eccf0;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb6acb030;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h25b5295a;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h62450461;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h6b0562a6;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h16a5ebdd;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'he1cf3ef7;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h1c599552;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hb057c849;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h555555fb;
          txc <= 4'h1;
          @ clk_0;
          txd <= 32'hd5555555;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h054e7c5f;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h0000588e;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hffffff00;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h8d2d0081;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h10000888;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h4dd00300;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00fe0000;
          txc <= 4'h4;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h00000000;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'hcb9286c3;
          txc <= 4'h0;
          @ clk_0;
          txd <= 32'h070707fd;
          txc <= 4'hf;
          @ clk_0;
        end

        txd <=32'h07070707;
        txc <=4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        if(EEE_ENABLED==1)
        begin
        txd <= 32'h0300009c;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'h0300009c;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'h0300009c;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'h0300009c;
        txc <= 4'h1;
        @ clk_0;
        end
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020103;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdbf64a6a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        if(EEE_ENABLED)
        begin
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h06060606;
          txc <= 4'hf;
          @ clk_0;
          txd <= 32'h07070707;
          txc <= 4'hf;
          @ clk_0;
        end
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h90642a00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7979deb6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h50ffef63;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc8b77608;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0038cc4d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7550843c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7d71c114;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcac14dc5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0fec8bb7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4208918d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'had8ecb72;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he6b68426;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020103;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h846e2e00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8f1a76c5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcd16bcd3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc2b3625f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h45446474;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8287c085;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h524f0a06;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5ceea67a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8b1bd5d5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf1775e7a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hda8ba833;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h24cb4ca0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5062bcc5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        if(EEE_ENABLED ==1)
        begin
        txd <= 32'h0300009c;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'h0300009c;
        txc <= 4'h1;
        @ clk_0;
        end
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020103;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6b972f00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcc9c9073;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfa0955db;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf4b5fe36;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h77a10621;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0976c772;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3e34469d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2d1ce9b4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2eb49825;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h04cdd9be;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha9d8287e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd1593bb9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0a298b6e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0707fd67;
        txc <= 4'he;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hccf13000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he6817350;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9d7247e2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hde6165fe;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha85cac50;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h48385d4c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf3cfd587;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf7dc6b7b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h08296d6e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb258fd3c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4f1e904c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hee5b753b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbe2d3d49;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h07fd36c6;
        txc <= 4'hc;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020103;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8c223100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9beabe2b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3342933e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9eaff703;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7a64b987;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8bbbed23;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h196ec3d2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd2d4b21d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hec5c4d73;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1733e274;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc9e0da2a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h87b6ba16;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd0f13f07;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfd22bbbd;
        txc <= 4'h8;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfb39dc05;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0c02ece6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbe85d57e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf3c87ea2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc877a5b1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3edbbaa2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hab482654;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc5a72762;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hddd40188;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdd10addc;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5f5df3ec;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h873e2731;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h13b81e0d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h846b0024;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf17b0c56;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hda8ac68b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0143b413;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h98ba271e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5d858a45;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h35e35f49;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h62bccda7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h49913070;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1c2b5c05;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2c1d81a6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbf214295;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6eee39b8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h76001118;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h152d441e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3f27de43;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5812f181;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4b3b4e76;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h82deeba2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h556627b7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4f7a478d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h036c85d0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4ae2eeea;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8805a91c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdf27e291;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h35ca964d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h33e077b3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha6ed4df0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1b381bfb;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h086b2a48;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h19c51f76;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h23a0ec62;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h25c32367;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h73179574;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd4e3c5cd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6d59f6fe;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4efb01cc;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h968a7bd3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd8b54542;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9af625c5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h078544ff;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h07b34611;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha6a9ab3a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h49cc153f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha4bf4f8a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4705c1c5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbf0137d5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h30ee1956;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0f64869b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcb80900b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h748067a3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8b1c2df6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4ada91a7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h099bac25;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1738bf8c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h50e3a556;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcc1e2e0a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h22c5c7ae;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h74068b03;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h83dccfb6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h37ce4425;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7fba79cf;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf0f999f5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbd4f74dc;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h608c2249;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h04c34fa8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5d6d2994;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6b0e52bf;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6e61c97e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4479e9e1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h55176889;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h272e19ef;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfa690a7a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4af342a6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'haeec0338;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7954f3d5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h11f5c6ef;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha7c37f23;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb7260de0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd672adf1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h353831cf;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc36e063b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf583b505;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5ef7fee5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc0837487;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h655ea9fb;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbd0c4cf4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3d15a249;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he31e2bcb;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc2b3c647;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h10c52d01;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9c799b0b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb44d74d0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h53d28556;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'haa0525a1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h92fa4e6a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03722718;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7266c34f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8ea0655f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf7e1320d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0af9b074;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4d00f46f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1db8619e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3d1796d0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h28939f6e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf10004e4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h93af8032;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha202e9f9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h227ceb82;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h05258d26;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5eb766da;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h946af8a9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h388b6ff1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5096d9c8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h86d37ee2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb4a98f96;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5072108a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2c71b01a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbb36ae4a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h208a7614;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6c9b0a23;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h97e39712;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd0d82fe1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5e0fc9f7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h90069b51;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb13930c3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h04e2a795;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha524a21f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hccf0a161;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3321b7f9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9656201f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6ec6282f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6a199236;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h80fad915;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h63f43d6d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h77337f9f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h89527a86;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc94c9b71;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9c0c04d2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h59bb7697;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6b5fe270;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf855fad3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h918695ce;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb6b91db8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h88e7cb53;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd886004d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h02c36d96;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcbff5967;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb148565e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h74deb082;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha52f1385;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf270dc0f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc4f455c2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5344ca7b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7636da72;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf35461dd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha5e69497;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h16164d90;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h817e49eb;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8dd5c242;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h894ee137;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h33f1534d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc22f9064;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h500f7dea;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1f3e46e5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbe3d2221;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4d9dab2a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdd71a582;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7fa32586;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'heffee072;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h65b270fd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3275be3d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h625f1b0e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0f1ceb0a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h83504901;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc4f27fc5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h59d8beb4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'heb0865a8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8a744904;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h312d45f3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he14bd994;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfeeed00c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h94ee68fc;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h53d0df58;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h93c50d72;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h27c5e108;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf9cfbe12;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8145c540;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb421b167;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbcd1a1b1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbf758aac;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hac886429;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h555b4771;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h40b3ca90;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he7715354;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc2731c44;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb5367831;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h71c9067b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6026ff70;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hafb4a027;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcb5f0c22;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd1744f8a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd35a7b0b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h85d13609;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h190c1403;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5f39e22d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h73449c08;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he8f85d47;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hde55362e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf580d090;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf0e7ea48;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcf4ad1d1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h060b1afd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h21f8c086;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7faa505b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd104ea9b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h93edfe77;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'had11a09b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'haeb4cf21;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h95719399;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf2f4d771;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h757c8163;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0b1c3082;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf4f5963f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8509b8bd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdb9f48e5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h037005de;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h84687850;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h02b15f6b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd8bf5065;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h55b310e0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2e5e9b7e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h134acff5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h73483ee1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h75c5c071;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6ee0ca51;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4ae68e27;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h847cb132;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hee6cd1e8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf6f56035;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfc70cf7f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3786c23b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4c979161;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha1c8f686;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb5e2fe21;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb55c5177;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h891090c6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h168b5764;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbc6c8261;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h537da5b0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2583957e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h14a177a6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfc281c0c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h05a1043a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h723c2fb7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdb673bdb;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd76c3dee;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he06fc619;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h42e2b0d9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h980c83c6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha2274b7e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbde69a8c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3556bad4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3aa8162b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h26845b01;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01bfe037;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h377011e7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3750a927;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd0679a53;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5ebee6f4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd3ca537c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h634d75c5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3f829566;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h155173b6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6dfee857;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h85a6f65e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hedcfef9e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8dcdb6ed;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5e0360ad;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7316150c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hde4dce64;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcd876b6b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3ffa4522;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd5c3d700;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfbc5ff41;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdf3ea6c3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h23115d7c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h12493f0b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h893cff05;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb4fcf11b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h65373c81;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9de6a179;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha25c3272;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h84667cca;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6acb8e13;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h439fcd41;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0bce6c81;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0e632174;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfbc7b13d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h99a2ccd8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h42b0681b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01362f7b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he99efcd2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd6e7236f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3bd1fb75;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2c1578a6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf00b1921;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3dfee41f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h05b6b707;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h28cba734;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf936df55;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfffc51f9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h89c5cdbf;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h20431fd7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h008ff387;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h660e9a95;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfdd8c74b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf2bb878d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb8cf29d4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h09930f07;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbcf0cb89;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h35297849;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hae32be8f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9bea699b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h09bf680d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h412fe3ca;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h35c90213;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha5ea3453;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb95fe55d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he5def62d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h56b935ee;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h872a8298;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1db21ff0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h741c7270;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2df14a51;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3e99d787;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hda952276;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfd63d201;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h632cac9f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h006cb1b4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc466f4ae;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h514b7faa;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he5c3e807;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc4fe82f4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd2656239;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6eefb2f1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8030ec4e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf1e04f85;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h64b42b2e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9de3da67;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc71df830;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hedbd896a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb29663d9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h63cb4c1a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h011c7994;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hae50d535;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd8dae25b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h015883ce;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h56b2f375;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha78b1f76;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h068d6598;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8273db2b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h67993302;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h07fdfda7;
        txc <= 4'hc;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020103;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdbf64a6a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020103;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5a1e0081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h336d292a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2b420081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb6d22a00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2754a7e6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb47d1985;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcc7f1cd5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5ccb1c41;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd52679ea;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3a56da3e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6521934b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h41f999ac;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf931e30b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4aff876b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h57eb499e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020103;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hccdb0081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3ab22e00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h53589720;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he63aaa7a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf6224983;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h781a6949;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h73a00bb1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8785f5e8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hea1f9c6d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h69452fe6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbfd72c53;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h99b1e338;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha5a41bed;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcea0c2b8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020103;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb3b50081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he4c72f00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha8403157;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9b9ed4d5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf361f5a6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfa91477e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc37b2ac3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2dcfe386;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcfd47d16;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h15b0fb1b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6924f823;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h99395b19;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h280447b4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6ae8b665;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0707fd55;
        txc <= 4'he;

        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020103;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb3b50081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he4c72f00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha8403157;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9b9ed4d5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf361f5a6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfa91477e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc37b2ac3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2dcfe386;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcfd47d16;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h15b0fb1b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6924f823;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h99395b19;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h280447b4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6ae8b665;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0707fd55;
        txc <= 4'he;


        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020103;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hde160081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb84a3000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0340bd22;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1ef5a243;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha931d85d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9f29a1ec;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8a260d2c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h83ea5e61;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc3765e0f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h68083d6d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfc5982f2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h640b8aa8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb47b21e1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha4f22e69;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h07fd78c8;
        txc <= 4'hc;
        
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020103;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hde160081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb84a3000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0340bd22;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1ef5a243;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha931d85d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9f29a1ec;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8a260d2c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h83ea5e61;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc3765e0f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h68083d6d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfc5982f2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h640b8aa8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb47b21e1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha4f22e69;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h07fd78c8;
        txc <= 4'hc;

@ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf4470081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h71533100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0484ff24;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2db50645;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h17c843dd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3ae122dd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h433f7438;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h245fe228;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8e04c4be;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4c366348;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h51f004fd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h19669700;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9a76d642;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6985b8cc;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfd873e82;
        txc <= 4'h8;

        
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf4470081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h71533100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0484ff24;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2db50645;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h17c843dd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3ae122dd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h433f7438;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h245fe228;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8e04c4be;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4c366348;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h51f004fd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h19669700;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9a76d642;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6985b8cc;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfd873e82;
        txc <= 4'h8;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03020100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000504;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h951d0081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h37fbdc05;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'haf764cca;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7d10a239;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h16c6f1fa;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h64d11226;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h34b1e35f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h041cbea5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h94fe707b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h92ebfb41;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h949cbe98;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf29587af;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbde7215c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf5ea4e5f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbdb47ff3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbb90e6b3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h35293c42;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h663c891e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha3c5940d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h09d26d97;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h33987bcc;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h41ef3ea7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8a3f8c6e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h323a5916;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7ad69306;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf3c629d3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01eee3b0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdcc72377;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h16ec169a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h47a1034d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdc43c29a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h17b4dff5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03a40e4a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6af685bb;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he8866fe1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha4b91511;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h52e3e95b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb752d311;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h34a14069;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1c3fdfba;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0e714b1d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3cb84e6f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h43afd084;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h918b810a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2bafceb3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3b4afe44;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h751ea682;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6d068782;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0680849d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4ec76955;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h52ce0c90;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h866d4cbd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h705847e7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h324e3b06;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'haa04d486;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb1411c4b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1c721828;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf2970839;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcb04d288;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4c462fe9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5da5efa9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5ca9453b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h581624d0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he3c94100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hda231b13;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4693d2b1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h16affb7d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h818b81b0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdc678a0e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'had3d272c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5251bbc5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h32f3bb07;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9bfcd3b3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h679d04e5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h67577a13;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'haaae0141;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc89d15cc;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h60546e21;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h75c9fa30;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8328c612;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h41e2ad14;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3bd83fde;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hddf0892a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbfae4408;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h82afd18b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5f748d6a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4c3d7e1a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h07f1a939;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3c4ce814;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hef24c176;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he4ab6317;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb204bc7b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3ec7b8ed;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8ce43ff6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0ba8677a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbe4db8ad;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hef898028;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcabf293a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5eca5d57;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h27cb5c93;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb43c7eba;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha2e037de;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hae712c3a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfa1f0eb1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0aae36b5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1dd0e9fd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3c0c01c6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h860983d5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6caae971;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbcf3ba59;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6db02dbc;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h40e75919;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hed03b0ef;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h52349b38;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdf6d1480;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h747f735c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1657e296;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h72586c33;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hef58c3fa;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hede8efe4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hdf4b4fc5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha3882411;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h11945444;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha841849a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7910361c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h62e978c7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha9343c58;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h89d8ba59;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf1771747;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h154f9368;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h40e44d34;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h05ce6b89;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h698eecb2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4a85f23c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3f5c1796;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb6756e38;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2cf6dcaa;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he98f97e0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h75eb72f2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hee078ec3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h18b82680;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h557d00a7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha091d4a1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he75583ff;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h63a155f8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3da3d463;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hacd06751;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3b07c2ce;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h19de5b32;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbabd0d4f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2d33e10e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h93e58ad6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc12edf9d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h67d425f2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h922d135f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd79215b6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h45169cbf;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h879d00eb;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h398c5d00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbaf30844;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1161b9c7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2719587d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hecd193e6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha1ff6be5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h95446e0f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbace7532;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb139183f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'haace58f9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf7e0eb27;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9039a8c9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf03355a2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7d87f110;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h348f45a6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc5fc2a48;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb5a75ab4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h445b30a6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha26ea238;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h64cfa359;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9df1a924;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h179e1d4b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0882c5b2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6e346b2d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb79c91c7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'haacf2547;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7aa33ede;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfd15e4ff;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h40b72db3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hefca8441;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4b0a8fd0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd91cc421;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1fab7322;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc8d1a7c1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h43211786;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4dee5ae1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7e05be9f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0b011884;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcc2cd72c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he1eea9a6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h11537d1e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1556d2a1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0219d4f5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9018be56;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hec9f24bd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf2476c08;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd9b8380f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8f5e47e5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbe81cd27;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h772668be;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf010b3f3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7ba89ea1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc58b9cae;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc8e7734f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc9de688a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb1d2c023;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7baff16a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h93a9b51b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h04b8de5a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1848a19f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h140d1680;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'haf163d18;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h69305934;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he68c61aa;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9cf13a16;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc4578fe4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h35a9ca88;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfec2ca9b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hde2533f7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h99de7f94;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h080bfff6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0c4de1cf;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha5fcff8c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h741c8187;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbefe3eea;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5dd0781b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha92bd3ce;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfea5807a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfa4de3b6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc1b5ae87;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h84f2b78b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3eac2dd4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h82c4d6e5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h400b0e86;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h977589c5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'haefc4558;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7ad5bd72;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6d2d4962;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5884fbc2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4424b276;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h62c73fce;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb16782df;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1283fd5d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h53c419bd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h89381540;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h163f1d38;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0fd1bae1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7c1dcb50;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd55e121d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h98619799;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9e2a7663;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h450e3555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h631cf688;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hba4e73b2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc6c7d5d1;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h173da3f6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc1f72f7f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h483d8971;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hddc1dafc;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h71092152;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hecac53b7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcb00f52e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcf187d53;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd5c8bbb3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5bf8bebe;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcb2e5b84;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfc3ec266;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9a411f08;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h402237d2;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc3a5aaf6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0a4a3e39;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h65c6c552;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf4d1f111;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h20102b75;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8b3b2f07;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6888ed3f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4a0a0050;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8d061f85;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h92919987;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8c9fe106;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4625fcbd;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf74b1d54;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h546fe640;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h06e106e4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03b8faa9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4d8c19e8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5ff7600b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc7a5c4e5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha7fd072b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h950e5939;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb98dbd34;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7a661784;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h779b55ba;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb3084849;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'heff7b5ab;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h884220ad;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd27d9e74;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb8d16d4a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha726fd97;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'haab3aa30;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd0f7922c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h19ccd173;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2f3370d7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha552a68b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h04f06ff0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h03b41fc4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbb37d5ff;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h601c93bb;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h345b3988;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hf4cbc114;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h41c18fb5;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6f898404;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hbc67e5ac;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3402be05;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h98312edf;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h045592a6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7eff2684;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h28e110ee;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h104c307e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2c5de71a;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h16785a36;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1ef1c130;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd28107ea;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hef61da07;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6ce228d6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfe8eb0b4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h09ab4938;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc404b60c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3d5798c4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb546c38d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9b2a2ad8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcb566aad;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h131c939c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb8185692;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h42f2df8e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1afe2277;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfb62c3c4;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h72ef39b0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h13664d88;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h66673d5d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4318f3d9;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h13f212ed;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h85f04569;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he3ffaca0;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0b4fb7ab;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h531081e8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h26632899;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h4d9df655;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3cb93139;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h0731c93b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd66d49b6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5a408cca;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'ha4ecf38f;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2564b00e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2edce969;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb9d4b339;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7a64f451;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'he045daac;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h10e51381;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2480dabf;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h58753de8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h3469325d;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h96b02d44;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h5f5a02d7;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h37208f30;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h276ae2e6;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2ccb5f83;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h7781b885;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8855f802;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h07fdd37e;
        txc <= 4'hc;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6a840081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2f6ef523;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcf7e0081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc35aad0b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9f210081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h55df1cc8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h459f0081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfd4da37c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9a960081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb1549d42;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6bc30081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfbc5491c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb2e20081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8419277e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h582b61e3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd60c8c15;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h582b61e3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1f389718;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd60c8c15;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h582b61e3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1f389718;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;       // end
        txc <= 4'hf;

        // Fault Sequences
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        
        // Added
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6a840081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2f6ef523;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcf7e0081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc35aad0b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9f210081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h55df1cc8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h459f0081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfd4da37c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9a960081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb1549d42;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6bc30081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfbc5491c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb2e20081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8419277e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h582b61e3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd60c8c15;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h582b61e3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000400;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9f15bc4e; // changed here
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000600;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h113251b8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h582b61e3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1f389718;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;   // end
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;

        // Added
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6a840081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h2f6ef523;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hcf7e0081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hc35aad0b;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9f210081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h55df1cc8;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h459f0081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfd4da37c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h9a960081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb1549d42;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h6bc30081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hfbc5491c;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hb2e20081;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h8419277e;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h582b61e3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd60c8c15;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h582b61e3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1f389718;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000200;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hd60c8c15;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h582b61e3;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h555555fb;
        txc <= 4'h1;
        @ clk_0;
        txd <= 32'hd5555555;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00c28001;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'hffffff00;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h01000888;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000100;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h00000000;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h1f389718;
        txc <= 4'h0;
        @ clk_0;
        txd <= 32'h070707fd;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;   // end

        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;

        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        
        

        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
        @ clk_0;
        txd <= 32'h07070707;
        txc <= 4'hf;
     end // initial begin
endmodule
