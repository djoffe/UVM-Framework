
import uvm_pkg::*;
import qvip_ahb_example_test_pkg::*;

module hvl_top;


initial run_test();

endmodule

